----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:16:46 11/16/2021 
-- Design Name: 
-- Module Name:    LUT6_beh - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LUT6_beh is
	GENERIC (
		INIT: STD_LOGIC_VECTOR (63 downto 0) := x"FF0000FFFF0000FF"
	);
   Port ( addr : in  STD_LOGIC_VECTOR (5 downto 0);
           Q : out  STD_LOGIC);
end LUT6_beh;

architecture Behavioral of LUT6_beh is
begin
	Q <= INIT(CONV_INTEGER(addr));
end Behavioral;

